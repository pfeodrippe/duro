module nao(x, z);
   input x;
   output z;

   assign z = x + 1;
endmodule
